`timescale 1ns / 1ps
//`include "user_module_341446083683025490.v"

module user_module_341446083683025490_tb;

    wire [7:0] io_in;
    wire [7:0] io_out;

    

endmodule
